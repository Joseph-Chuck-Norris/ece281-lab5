--+----------------------------------------------------------------------------
--|
--| NAMING CONVENSIONS :
--|
--|    xb_<port name>           = off-chip bidirectional port ( _pads file )
--|    xi_<port name>           = off-chip input port         ( _pads file )
--|    xo_<port name>           = off-chip output port        ( _pads file )
--|    b_<port name>            = on-chip bidirectional port
--|    i_<port name>            = on-chip input port
--|    o_<port name>            = on-chip output port
--|    c_<signal name>          = combinatorial signal
--|    f_<signal name>          = synchronous signal
--|    ff_<signal name>         = pipeline stage (ff_, fff_, etc.)
--|    <signal name>_n          = active low signal
--|    w_<signal name>          = top level wiring signal
--|    g_<generic name>         = generic
--|    k_<constant name>        = constant
--|    v_<variable name>        = variable
--|    sm_<state machine type>  = state machine type definition
--|    s_<signal name>          = state name
--|
--+----------------------------------------------------------------------------
--|
--| ALU OPCODES:
--|
--|     ADD     000
--|
--|
--|
--|
--+----------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;


entity ALU is
    port (
    i_A : in STD_LOGIC_VECTOR (7 DOWNTO 0);
    i_B : in STD_LOGIC_VECTOR (7 DOWNTO 0);
    i_op : in STD_LOGIC_VECTOR (2 DOWNTO 0);
    o_results : out STD_LOGIC_VECTOR (7 DOWNTO 0);
    o_flags : out STD_LOGIC_VECTOR (2 DOWNTO 0)
    );
end ALU;

architecture behavioral of ALU is 
  
	-- declare components and signals
    signal w_decoderOne : STD_LOGIC_VECTOR(7 DOWNTO 0);
    signal w_adder : STD_LOGIC_VECTOR(7 DOWNTO 0);
    signal w_SEL : STD_LOGIC_VECTOR(1 DOWNTO 0);
    signal w_D_IN : STD_LOGIC_VECTOR(3 DOWNTO 0);

    
begin
	-- PORT MAPS ----------------------------------------
	    w_decoderOne <= not i_B when i_op(2) = '1' else 
	                 i_B;
        w_adder <= (i_A XOR w_decoderOne) OR i_op(2);
        
        with w_SEL select
            o_results <= w_adder when "00",
--                          when "01",
--                          when "10",
--                          when "11",
                         "00000000" when others;
	
	
	-- CONCURRENT STATEMENTS ----------------------------
	   o_flags[0] <= i_results(7);
	   o_flags[1] <= not (i_results or i_results);
	   
	
	
end behavioral;
